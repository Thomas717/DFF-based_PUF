VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM256
  CLASS BLOCK ;
  FOREIGN RAM256 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1971.200 BY 799.680 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.452000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 85.120 1971.200 85.680 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.452000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 142.240 1971.200 142.800 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.452000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 199.360 1971.200 199.920 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.452000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 256.480 1971.200 257.040 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.452000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 313.600 1971.200 314.160 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.452000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 370.720 1971.200 371.280 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.452000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 427.840 1971.200 428.400 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.132000 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 484.960 1971.200 485.520 ;
    END
  END A0[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.366000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 542.080 1971.200 542.640 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 646.240 0.000 646.800 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 707.840 0.000 708.400 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 769.440 0.000 770.000 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 831.040 0.000 831.600 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 892.640 0.000 893.200 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 954.240 0.000 954.800 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1015.840 0.000 1016.400 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1077.440 0.000 1078.000 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1139.040 0.000 1139.600 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1200.640 0.000 1201.200 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 0.000 92.400 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1262.240 0.000 1262.800 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1323.840 0.000 1324.400 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1385.440 0.000 1386.000 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1447.040 0.000 1447.600 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1508.640 0.000 1509.200 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1570.240 0.000 1570.800 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1631.840 0.000 1632.400 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1693.440 0.000 1694.000 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1755.040 0.000 1755.600 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1816.640 0.000 1817.200 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 0.000 154.000 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1878.240 0.000 1878.800 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1939.840 0.000 1940.400 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 0.000 215.600 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 0.000 277.200 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 0.000 338.800 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 0.000 400.400 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 461.440 0.000 462.000 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 523.040 0.000 523.600 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 0.000 585.200 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 797.680 30.800 799.680 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 646.240 797.680 646.800 799.680 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 707.840 797.680 708.400 799.680 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 769.440 797.680 770.000 799.680 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 831.040 797.680 831.600 799.680 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 892.640 797.680 893.200 799.680 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 954.240 797.680 954.800 799.680 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1015.840 797.680 1016.400 799.680 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1077.440 797.680 1078.000 799.680 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1139.040 797.680 1139.600 799.680 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1200.640 797.680 1201.200 799.680 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 797.680 92.400 799.680 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1262.240 797.680 1262.800 799.680 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1323.840 797.680 1324.400 799.680 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1385.440 797.680 1386.000 799.680 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1447.040 797.680 1447.600 799.680 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1508.640 797.680 1509.200 799.680 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1570.240 797.680 1570.800 799.680 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1631.840 797.680 1632.400 799.680 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1693.440 797.680 1694.000 799.680 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1755.040 797.680 1755.600 799.680 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1816.640 797.680 1817.200 799.680 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 797.680 154.000 799.680 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1878.240 797.680 1878.800 799.680 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1939.840 797.680 1940.400 799.680 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 797.680 215.600 799.680 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 797.680 277.200 799.680 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 797.680 338.800 799.680 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 797.680 400.400 799.680 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 461.440 797.680 462.000 799.680 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 523.040 797.680 523.600 799.680 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 797.680 585.200 799.680 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.048000 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 28.000 1971.200 28.560 ;
    END
  END EN0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.320 3.620 19.920 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 171.920 3.620 173.520 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 325.520 3.620 327.120 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 479.120 3.620 480.720 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 632.720 3.620 634.320 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 786.320 3.620 787.920 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 939.920 3.620 941.520 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1093.520 3.620 1095.120 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1247.120 3.620 1248.720 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1400.720 3.620 1402.320 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1554.320 3.620 1555.920 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1707.920 3.620 1709.520 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1861.520 3.620 1863.120 796.060 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 95.120 3.620 96.720 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 248.720 3.620 250.320 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 402.320 3.620 403.920 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 555.920 3.620 557.520 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 709.520 3.620 711.120 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 863.120 3.620 864.720 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1016.720 3.620 1018.320 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1170.320 3.620 1171.920 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1323.920 3.620 1325.520 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1477.520 3.620 1479.120 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1631.120 3.620 1632.720 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1784.720 3.620 1786.320 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1938.320 3.620 1939.920 796.060 ;
    END
  END VSS
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.452000 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 599.200 1971.200 599.760 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.452000 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 656.320 1971.200 656.880 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.452000 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 713.440 1971.200 714.000 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.452000 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.200 770.560 1971.200 771.120 ;
    END
  END WE0[3]
  OBS
      LAYER Metal1 ;
        RECT 2.800 3.620 1968.400 796.060 ;
      LAYER Metal2 ;
        RECT 0.700 797.380 29.940 799.590 ;
        RECT 31.100 797.380 91.540 799.590 ;
        RECT 92.700 797.380 153.140 799.590 ;
        RECT 154.300 797.380 214.740 799.590 ;
        RECT 215.900 797.380 276.340 799.590 ;
        RECT 277.500 797.380 337.940 799.590 ;
        RECT 339.100 797.380 399.540 799.590 ;
        RECT 400.700 797.380 461.140 799.590 ;
        RECT 462.300 797.380 522.740 799.590 ;
        RECT 523.900 797.380 584.340 799.590 ;
        RECT 585.500 797.380 645.940 799.590 ;
        RECT 647.100 797.380 707.540 799.590 ;
        RECT 708.700 797.380 769.140 799.590 ;
        RECT 770.300 797.380 830.740 799.590 ;
        RECT 831.900 797.380 892.340 799.590 ;
        RECT 893.500 797.380 953.940 799.590 ;
        RECT 955.100 797.380 1015.540 799.590 ;
        RECT 1016.700 797.380 1077.140 799.590 ;
        RECT 1078.300 797.380 1138.740 799.590 ;
        RECT 1139.900 797.380 1200.340 799.590 ;
        RECT 1201.500 797.380 1261.940 799.590 ;
        RECT 1263.100 797.380 1323.540 799.590 ;
        RECT 1324.700 797.380 1385.140 799.590 ;
        RECT 1386.300 797.380 1446.740 799.590 ;
        RECT 1447.900 797.380 1508.340 799.590 ;
        RECT 1509.500 797.380 1569.940 799.590 ;
        RECT 1571.100 797.380 1631.540 799.590 ;
        RECT 1632.700 797.380 1693.140 799.590 ;
        RECT 1694.300 797.380 1754.740 799.590 ;
        RECT 1755.900 797.380 1816.340 799.590 ;
        RECT 1817.500 797.380 1877.940 799.590 ;
        RECT 1879.100 797.380 1939.540 799.590 ;
        RECT 1940.700 797.380 1971.060 799.590 ;
        RECT 0.700 2.300 1971.060 797.380 ;
        RECT 0.700 0.090 29.940 2.300 ;
        RECT 31.100 0.090 91.540 2.300 ;
        RECT 92.700 0.090 153.140 2.300 ;
        RECT 154.300 0.090 214.740 2.300 ;
        RECT 215.900 0.090 276.340 2.300 ;
        RECT 277.500 0.090 337.940 2.300 ;
        RECT 339.100 0.090 399.540 2.300 ;
        RECT 400.700 0.090 461.140 2.300 ;
        RECT 462.300 0.090 522.740 2.300 ;
        RECT 523.900 0.090 584.340 2.300 ;
        RECT 585.500 0.090 645.940 2.300 ;
        RECT 647.100 0.090 707.540 2.300 ;
        RECT 708.700 0.090 769.140 2.300 ;
        RECT 770.300 0.090 830.740 2.300 ;
        RECT 831.900 0.090 892.340 2.300 ;
        RECT 893.500 0.090 953.940 2.300 ;
        RECT 955.100 0.090 1015.540 2.300 ;
        RECT 1016.700 0.090 1077.140 2.300 ;
        RECT 1078.300 0.090 1138.740 2.300 ;
        RECT 1139.900 0.090 1200.340 2.300 ;
        RECT 1201.500 0.090 1261.940 2.300 ;
        RECT 1263.100 0.090 1323.540 2.300 ;
        RECT 1324.700 0.090 1385.140 2.300 ;
        RECT 1386.300 0.090 1446.740 2.300 ;
        RECT 1447.900 0.090 1508.340 2.300 ;
        RECT 1509.500 0.090 1569.940 2.300 ;
        RECT 1571.100 0.090 1631.540 2.300 ;
        RECT 1632.700 0.090 1693.140 2.300 ;
        RECT 1694.300 0.090 1754.740 2.300 ;
        RECT 1755.900 0.090 1816.340 2.300 ;
        RECT 1817.500 0.090 1877.940 2.300 ;
        RECT 1879.100 0.090 1939.540 2.300 ;
        RECT 1940.700 0.090 1971.060 2.300 ;
      LAYER Metal3 ;
        RECT 0.650 771.420 1971.110 799.540 ;
        RECT 0.650 770.260 1968.900 771.420 ;
        RECT 0.650 714.300 1971.110 770.260 ;
        RECT 0.650 713.140 1968.900 714.300 ;
        RECT 0.650 657.180 1971.110 713.140 ;
        RECT 0.650 656.020 1968.900 657.180 ;
        RECT 0.650 600.060 1971.110 656.020 ;
        RECT 0.650 598.900 1968.900 600.060 ;
        RECT 0.650 542.940 1971.110 598.900 ;
        RECT 0.650 541.780 1968.900 542.940 ;
        RECT 0.650 485.820 1971.110 541.780 ;
        RECT 0.650 484.660 1968.900 485.820 ;
        RECT 0.650 428.700 1971.110 484.660 ;
        RECT 0.650 427.540 1968.900 428.700 ;
        RECT 0.650 371.580 1971.110 427.540 ;
        RECT 0.650 370.420 1968.900 371.580 ;
        RECT 0.650 314.460 1971.110 370.420 ;
        RECT 0.650 313.300 1968.900 314.460 ;
        RECT 0.650 257.340 1971.110 313.300 ;
        RECT 0.650 256.180 1968.900 257.340 ;
        RECT 0.650 200.220 1971.110 256.180 ;
        RECT 0.650 199.060 1968.900 200.220 ;
        RECT 0.650 143.100 1971.110 199.060 ;
        RECT 0.650 141.940 1968.900 143.100 ;
        RECT 0.650 85.980 1971.110 141.940 ;
        RECT 0.650 84.820 1968.900 85.980 ;
        RECT 0.650 28.860 1971.110 84.820 ;
        RECT 0.650 27.700 1968.900 28.860 ;
        RECT 0.650 0.140 1971.110 27.700 ;
      LAYER Metal4 ;
        RECT 5.180 796.360 1965.460 799.590 ;
        RECT 5.180 3.320 18.020 796.360 ;
        RECT 20.220 3.320 94.820 796.360 ;
        RECT 97.020 3.320 171.620 796.360 ;
        RECT 173.820 3.320 248.420 796.360 ;
        RECT 250.620 3.320 325.220 796.360 ;
        RECT 327.420 3.320 402.020 796.360 ;
        RECT 404.220 3.320 478.820 796.360 ;
        RECT 481.020 3.320 555.620 796.360 ;
        RECT 557.820 3.320 632.420 796.360 ;
        RECT 634.620 3.320 709.220 796.360 ;
        RECT 711.420 3.320 786.020 796.360 ;
        RECT 788.220 3.320 862.820 796.360 ;
        RECT 865.020 3.320 939.620 796.360 ;
        RECT 941.820 3.320 1016.420 796.360 ;
        RECT 1018.620 3.320 1093.220 796.360 ;
        RECT 1095.420 3.320 1170.020 796.360 ;
        RECT 1172.220 3.320 1246.820 796.360 ;
        RECT 1249.020 3.320 1323.620 796.360 ;
        RECT 1325.820 3.320 1400.420 796.360 ;
        RECT 1402.620 3.320 1477.220 796.360 ;
        RECT 1479.420 3.320 1554.020 796.360 ;
        RECT 1556.220 3.320 1630.820 796.360 ;
        RECT 1633.020 3.320 1707.620 796.360 ;
        RECT 1709.820 3.320 1784.420 796.360 ;
        RECT 1786.620 3.320 1861.220 796.360 ;
        RECT 1863.420 3.320 1938.020 796.360 ;
        RECT 1940.220 3.320 1965.460 796.360 ;
        RECT 5.180 0.090 1965.460 3.320 ;
  END
END RAM256
END LIBRARY

